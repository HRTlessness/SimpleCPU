module control(input clk, input reset);

endmodule
